-- Part of TDT4255 Computer Design laboratory exercises
-- Group for Computer Architecture and Design
-- Department of Computer and Information Science
-- Norwegian University of Science and Technology

-- MIPSProcessor.vhd
-- The MIPS processor component to be used in Exercise 1 and 2.

-- TODO replace the architecture DummyArch with a working Behavioral

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity MIPSProcessor is
	generic (
		ADDR_WIDTH 		: integer := 8;
		ADDR_REG_WIDTH : integer := 5;
		DATA_WIDTH 		: integer := 32;
		regfile_size 	: natural := 32);
	port ( 
		clk, reset 				: in std_logic;
		processor_enable		: in std_logic;
		imem_data_in			: in std_logic_vector(DATA_WIDTH-1 downto 0);
		imem_address			: out std_logic_vector(ADDR_WIDTH-1 downto 0);
		dmem_data_in			: in std_logic_vector(DATA_WIDTH-1 downto 0);
		dmem_address			: out std_logic_vector(ADDR_WIDTH-1 downto 0);
		dmem_data_out			: out std_logic_vector(DATA_WIDTH-1 downto 0);
		dmem_write_enable		: out std_logic
	);
end MIPSProcessor;

architecture Behavioral of MIPSProcessor is
	
	-- PC signals
	signal address_in		: std_logic_vector(DATA_WIDTH-1 downto 0);
	signal address_out	: std_logic_vector(DATA_WIDTH-1 downto 0);
	signal next_address  : std_logic_vector(DATA_WIDTH-1 downto 0);
	--ALU PC  signal
	signal empty : boolean;
	-- IF_ID_Register 
	signal instruction : std_logic_vector(DATA_WIDTH-1 downto 0);
	signal pc_address : std_logic_vector(DATA_WIDTH-1 downto 0);
	-- registers signals
	signal read_data_1	: std_logic_vector(DATA_WIDTH-1 downto 0);
	signal read_data_2	: std_logic_vector(DATA_WIDTH-1 downto 0);
	signal write_data    : std_logic_vector(DATA_WIDTH-1 downto 0);
   signal write_reg_add :  std_logic_vector(ADDR_REG_WIDTH-1 downto 0);	
	-- ID_EX_Register
	signal pc_address_ex  : std_logic_vector(31 downto 0);
	signal read_data_1_ex : std_logic_vector(31 downto 0);
	signal read_data_2_ex : std_logic_vector(31 downto 0);
	signal extended_value_ex : std_logic_vector(31 downto 0);
	signal instruction_20to16_ex : std_logic_vector(4 downto 0);
	signal instruction_15to11_ex : std_logic_vector(4 downto 0);
	-- EX_MEM_Register
	signal add_result : std_logic_vector(DATA_WIDTH-1 downto 0);
	signal zero_out : std_logic;
	signal alu_result_mem : std_logic_vector(31 downto 0);
	signal write_register_mem : std_logic_vector(31 downto 0);
	signal reg_write_mem : std_logic;
   signal branch_mem : std_logic;
   

	-- control signal outputs
	signal regwrite_ex : STD_LOGIC;
	signal branch_ex	 : STD_LOGIC;
	signal regdst_ex	 : STD_LOGIC;
	signal aluop_ex	 : std_logic_vector(1 downto 0);
	signal alusrc_ex	 : STD_LOGIC;
	signal memwrite_ex : STD_LOGIC;
	signal memtoreg_ex : STD_LOGIC;
	-- ALU signals
	signal zero			: boolean;	
	signal data_2     : std_logic_vector(DATA_WIDTH-1 downto 0);
	signal alu_result : std_logic_vector(DATA_WIDTH-1 downto 0); -- BECAREFUL alu result is a buffer signal
	-- ALU Control signal
	signal alu_op     : std_logic_vector(3 downto 0); 
	-- Control unit signals
	signal reg_write  : std_logic :='0';
	signal op_code    : std_logic_vector(1 downto 0):="00";
	signal reg_dst    : std_logic :='0';
	signal branch     : std_logic :='0';
	signal jump			: std_logic :='0';
	signal mem_to_reg : std_logic :='0';
	signal alu_src    : std_logic :='0';
	-- SignExtend
	signal extend_out : std_logic_vector(DATA_WIDTH-1 downto 0);
	
	
begin
	
	-- Mux before Program counter
	
	
	
	add_result <= 	std_logic_vector(signed(pc_address_ex) + signed(extended_value_ex));				
	-- Mux before regfile
	write_reg_add <=	instruction_20to16_ex when regdst_ex='0' else
							instruction_15to11_ex; 
	-- Mux before ALU
	data_2 <= 	read_data_2_ex when alusrc_ex='0' else
					extended_value_ex; 
	-- Mux after Data memory
	write_data <= 	alu_result when mem_to_reg='0' else 
						dmem_data_in; 
						
	imem_address <= address_out(ADDR_WIDTH-1 downto 0);
	dmem_address <= alu_result(ADDR_WIDTH-1 downto 0);
	dmem_data_out<= read_data_2;
	
	
	IF_ID_Register : entity work.if_id_reg 
	port map(
		clk						=> clk,
		rst						=> reset,
		imem_instruction_in	=> imem_data_in,
		pc_address_in			=> next_address,
		imem_instruction_out	=> instruction,
		pc_address_out			=> pc_address);
	
	ID_EX_Register : entity work.id_ex_reg
  	port map (
		-- inputs
      clk			   => clk,
		rst			   => reset,
		pc_address_in  => pc_address,
		read_data_1_in => read_data_1,
		read_data_2_in => read_data_2,
		extended_value_in => extend_out,
		instruction_20to16_in => instruction(20 downto 16),
		instruction_15to11_in => instruction(15 downto 11),
		
		--control signal inputs
		regwrite_in => reg_write,
		branch_in	=> branch,
		regdst_in	=> reg_dst,
		aluop_in	=> op_code,
		alusrc_in	=> alu_src,
		memwrite_in => mem_write,
		memtoreg_in => mem_to_reg,
		
		-- outputs
		pc_address_out  => pc_address_ex,
		read_data_1_out => read_data_1_ex,
		read_data_2_out => read_data_2_ex,
		extended_value_out => extended_value_ex,
		instruction_20to16_out =>instruction_20to16_ex,
		instruction_15to11_out => instruction_15to11_ex,
		
		-- control signal outputs
		regwrite_out => regwrite_ex,
		branch_out	 => branch_ex,
		regdst_out	 => regdst_ex,
		aluop_out	 => aluop_ex,
		alusrc_out	 => alusrc_ex,
		memwrite_out => memwrite_ex,
		memtoreg_out => memtoreg_ex,
		
    --for forwarding unit
    reg_rt_in => ,
    reg_rt_out => ,
    reg_rs_in => ,
    reg_rs_out => );
	
	 
	 EX_MEM_Register : entity work.ex_to_mem 
    port (
        clk  => clk,
        rst  => reset,
        add_result_in => add_result,
        add_result_out  => add_result_mem,
        zero_in  => zero, 
        zero_out => zero_mem,
        alu_result_in  => alu_result,
        alu_result_out => alu_result_mem,
        read_data_in  => read_data_2_ex,
        read_data_out => read_data_mem,
        write_register_in => write_reg_add,
        write_register_out => write_register_mem,

        --control
        reg_write_in  => regwrite_ex,
        reg_write_out  => dmem_data_out,
        branch_in  => branch_ex,
        branch_out => branch_mem,
        mem_to_reg_in  => memtoreg_ex,
        mem_to_reg_out => memtoreg_mem,   
        mem_write_in => memwrite_ex,
        mem_write_out => dmem_write_enable
    );
	 
	MEM_WB_Register : entity work.mem_to_wb
    port map(
        clk => clk,
        rst => reset,
        alu_result_in => read_data_mem,
        alu_result_out => ,
        write_register_in => write_register_mem,
        write_register_out => ,
		  mem_to_reg_in  => memtoreg_ex,
        mem_to_reg_out =>
    ); 
	 
	SignExtend : entity work.SignExtend
		port map( 
			data_in  => instruction( 15 downto 0),
         data_out => extend_out);
	
	RegisterFile : entity work.RegisterFile
		generic map(
			ADDR_REG_WIDTH => ADDR_REG_WIDTH,
			DATA_WIDTH => DATA_WIDTH,
			size => regfile_size )
		port map(
			clk => clk,
			rst	=> reset,
			RegWrite => reg_write,		
			read_register1_addr => instruction( 25 downto 21), 
			read_register2_addr => instruction( 20 downto 16),
			write_register_addr => write_reg_add,
			write_data	=> write_data,
			read_data1	=> read_data_1,
			read_data2	=> read_data_2);
		
	ALU : entity work.ALU
		port map (
			rt  			=> read_data_1_ex,
			rs				=> data_2,
			alu_op		=> alu_op ,
			alu_result	=> alu_result,
			zero			=> zero );
	
	ALU_PC : entity work.ALU
		port map (
			rt  			=> address_out,
			rs				=> x"00000001",
			alu_op		=> "0010" ,
			alu_result	=> next_address,
			zero			=> empty);
			
	ALU_Ctrl : entity work.ALU_Ctrl
		port map(
			op_code => aluop_ex,
			instruction_funct => instruction( 5 downto 0) ,			
			alu_op =>  alu_op);
	
	program_counter : entity work.program_counter
		port map(
			clk      => clk,
			rst		=> reset,
			write_en => write_en,	
			PC_in		=> address_in,
			PC_out	=> address_out); 	
			
	control_unit : entity work.control_unit
		port map(
		 clk => clk,
		 rst => reset,	  
		 instruction => instruction(31 downto 26),
		 reg_dst    => reg_dst,
		 branch     => branch,
		 jump			=> jump,
		 mem_to_reg  => mem_to_reg,
		 alu_op      => op_code ,
		 alu_src     => alu_src,
		 reg_write   => reg_write ,
		 mem_write   => dmem_write_enable,
		 processor_enable => processor_enable	);	
	
end Behavioral;

